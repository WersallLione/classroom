module mux2(
input wire FPGA_CLK    ,
input wire en_key      ,
input wire din1        ,
input wire din2,       ,

output reg [3:0] dout
);

endmodule